class or_sequence
