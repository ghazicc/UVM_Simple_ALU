class subtraction
